library verilog;
use verilog.vl_types.all;
entity hello_world_vlg_check_tst is
    port(
        Sand            : in     vl_logic;
        Sor             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end hello_world_vlg_check_tst;
