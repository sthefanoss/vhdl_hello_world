library verilog;
use verilog.vl_types.all;
entity hello_world_vlg_vec_tst is
end hello_world_vlg_vec_tst;
